module comparison_module (input1, input2, eq, gt, lt);
	input [2:0] input1;
	input [2:0] input2;
	output eq, gt, lt;

    assign eq = input1 == input2;
    assign gt = input1 > input2;
    assign lt = input1 < input2;

endmodule
