module ones_counter(
    input [3:0] in,
    output reg [3:0] count
);

	// * means if anythoing changes, called wildcard?
	always @(*) begin
		count = in[0] + in[1] + in[2] + in[3];
	end

endmodule