module sequence_detector_part_2 (SW, KEY, LEDR);
	// TODO: define input and output ports:
	input [1:0] SW;
   input [0:0] KEY;
   output [9:0] LEDR;
	// y_Q  current state, y_D  next state
	reg [3:0] y_Q, y_D;
	
   wire Clock, Resetn, w;
   reg out;

   assign Clock = ~KEY[0];
   assign Resetn = SW[0];
   assign w = SW[1];
	
	
	// define state parameters:
	parameter A = 4'b0000, B = 4'b0001, C = 4'b0010, D = 4'b0011, E = 4'b0100, F = 4'b0101, G = 4'b0110, H = 4'b0111, I = 4'b1000;
	
	// TODO: implement the state table:
		always @(w, y_Q) begin 
		case (y_Q)
			A: if (!w) y_D <= B; else y_D <= F;
			// for 000
			B: if (!w) y_D <= C; else y_D <= F;
         C: if (!w) y_D <= D; else y_D <= F;
         D: if (!w) y_D <= E; else y_D <= F;
         E: if (!w) y_D <= E; else y_D <= F;
			// for 111
         F: if (!w) y_D <= B; else y_D <= G;
         G: if (!w) y_D <= B; else y_D <= H;
         H: if (!w) y_D <= B; else y_D <= I;
         I: if (!w) y_D <= B; else y_D <= I;
			// idk if I need this but just in case
			default: y_D <= 4'bxxxx;
		endcase
	end

	// TODO: udpate the state on rising clock edges:
	always @(posedge Clock) begin: state_FFs
			if (Resetn)
				y_Q <= A;
			else
            y_Q <= y_D;
    end // state_FFS

    // output logic
    always @(y_Q) begin
        case (y_Q)
            E: out <= 1'b1;
				I: out <= 1'b1;
            default: out <= 1'b0;
        endcase
    end


	// TODO: assignments for output and the LEDs:
	 assign LEDR[3:0] = y_Q;
    assign LEDR[9] = out; 
	
endmodule